// Mohammad Abu Shams.
// All ciruits using a structural model.
module Circuit(A,B,C0,S,Cout);
input [3:0] B,A;
input C0;
output Cout;
output[3:0]S;
wire [3:0] I1,F;

Complement G1(B[3],B[2],B[1],B[0],I1[3],I1[2],I1[1],I1[0]);
QMUX G2(B,I1,C0,F);
BCDA G3(A,F,C0,S,Cout);
endmodule
